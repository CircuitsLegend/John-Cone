// This module uses behavioral Verilog.
//
// Behavior:
//    If "en" (enable) is 1, then input d is 
//    written to output q with a one-cycle delay.
//
//    If "en" is 0, then q is reset to 0 with
//    a one-cycle delay.
//      
//      `
`timescale 1ns/1ps
module simple_module (
		      input clk,
		      input en,
		      input d,
		      output reg q
		      );

   initial q=0;
   
   always @(posedge clk) begin
      if (en)
	q <= d;   // NON-BLOCKING ASSIGNMENT specifies D Flip Flop
      else        // The flip-flop creates a one-cycle delay before
	q <= q;   // q is changed
   end
endmodule // simple_module
