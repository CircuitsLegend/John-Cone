Use `include to include the reverse_bits_function in a top module called reverse_bits_module
Instead of task invocations, use the function syntax:
   q = reverse_bits_function(a);
